-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.1.0 Build 162 10/23/2013 SJ Web Edition"
-- CREATED		"Sun Sep 18 09:01:10 2022"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY mx2x8 IS 
	PORT
	(
		EN :  IN  STD_LOGIC;
		S0 :  IN  STD_LOGIC;
		I0 :  IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		I1 :  IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		Y :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END mx2x8;

ARCHITECTURE bdf_type OF mx2x8 IS 

SIGNAL	Y_ALTERA_SYNTHESIZED :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;


BEGIN 



SYNTHESIZED_WIRE_16 <= I0(0) AND EN AND SYNTHESIZED_WIRE_24;


SYNTHESIZED_WIRE_24 <= NOT(S0);



Y_ALTERA_SYNTHESIZED(7) <= SYNTHESIZED_WIRE_1 OR SYNTHESIZED_WIRE_2;


Y_ALTERA_SYNTHESIZED(6) <= SYNTHESIZED_WIRE_3 OR SYNTHESIZED_WIRE_4;


Y_ALTERA_SYNTHESIZED(5) <= SYNTHESIZED_WIRE_5 OR SYNTHESIZED_WIRE_6;


Y_ALTERA_SYNTHESIZED(4) <= SYNTHESIZED_WIRE_7 OR SYNTHESIZED_WIRE_8;


Y_ALTERA_SYNTHESIZED(3) <= SYNTHESIZED_WIRE_9 OR SYNTHESIZED_WIRE_10;


Y_ALTERA_SYNTHESIZED(2) <= SYNTHESIZED_WIRE_11 OR SYNTHESIZED_WIRE_12;


Y_ALTERA_SYNTHESIZED(1) <= SYNTHESIZED_WIRE_13 OR SYNTHESIZED_WIRE_14;


Y_ALTERA_SYNTHESIZED(0) <= SYNTHESIZED_WIRE_15 OR SYNTHESIZED_WIRE_16;


SYNTHESIZED_WIRE_14 <= I0(1) AND EN AND SYNTHESIZED_WIRE_24;


SYNTHESIZED_WIRE_12 <= I0(2) AND EN AND SYNTHESIZED_WIRE_24;


SYNTHESIZED_WIRE_10 <= I0(3) AND EN AND SYNTHESIZED_WIRE_24;


SYNTHESIZED_WIRE_8 <= I0(4) AND EN AND SYNTHESIZED_WIRE_24;


SYNTHESIZED_WIRE_6 <= I0(5) AND EN AND SYNTHESIZED_WIRE_24;


SYNTHESIZED_WIRE_4 <= I0(6) AND EN AND SYNTHESIZED_WIRE_24;


SYNTHESIZED_WIRE_2 <= I0(7) AND EN AND SYNTHESIZED_WIRE_24;


SYNTHESIZED_WIRE_15 <= I1(0) AND EN AND S0;


SYNTHESIZED_WIRE_13 <= I1(1) AND EN AND S0;


SYNTHESIZED_WIRE_11 <= I1(2) AND EN AND S0;


SYNTHESIZED_WIRE_9 <= I1(3) AND EN AND S0;


SYNTHESIZED_WIRE_7 <= I1(4) AND EN AND S0;


SYNTHESIZED_WIRE_5 <= I1(5) AND EN AND S0;


SYNTHESIZED_WIRE_3 <= I1(6) AND EN AND S0;


SYNTHESIZED_WIRE_1 <= I1(7) AND EN AND S0;

Y <= Y_ALTERA_SYNTHESIZED;

END bdf_type;